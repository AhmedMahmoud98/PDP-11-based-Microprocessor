LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

-- Control Store Data
ENTITY ROM IS
	PORT(   
                address : IN  std_logic_vector(4 DOWNTO 0);
		micro_instruction : OUT std_logic_vector(19 DOWNTO 0)
	    );
END ENTITY ROM;

ARCHITECTURE ROM_arch OF ROM IS
TYPE ROM_memory IS ARRAY ( 0 to 2**5 - 1) of std_logic_vector(19 downto 0);
  CONSTANT ROM_data : ROM_memory := (
    	0  => "11000010011010110000",
		1  => "01011110011010000000",
		2  => "01010110011111000111",
		3  => "00110110000010000000",
		4  => "10110110100011110011",
		5  => "00000000011001110011",
		6  => "00111110010110110011",
		7  => "01000110001011110011",
		8  => "01001110100111001011",
		9  => "11000001010010110000",
		10 => "11000001010010010000",
		11 => "11000001010111010011",
		12 => "10010110101111010011",
		13 => "01110110000011110011",
		14 => "01111110110111001011",
		15 => "10010110010110110011",
		16 => "10010110010111010011",
		17 => "10010110010100110001",
		18 => "10011110000010000000",
		19 => "10100110010110110011",
		20 => "00000101001101110011",
		21 => "00000000111111110010",
		22 => "10000100101111001111",
		23 => "00000111111111110011",
		24 => "10110110001011110011",
		25 => "11000011001010110000",
		26 => "10010110101100110001",
		27 => "11010110001010110011",
		28 => "00000000001001110011",
		29 => "00000111111111110011",
		30 => "00000111111111110011",
		31 => "11111110111111110011"
			);

BEGIN
	micro_instruction <= ROM_data(to_integer(unsigned(address)));
END ROM_arch;

